module tb_snow_vi_aes_round();
endmodule // tb_snow_vi_aes_round
