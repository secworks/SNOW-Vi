module tb_snow_vi_core();
endmodule // tb_snow_vi_core
