module tb_snow_vi();
endmodule // tb_snow_vi
